module calculator (
    input  logic       clk_i,
    input  logic       rst_i,

    input  logic [4:0] a_i,
    input  logic [4:0] b_i,
    input  logic       input_valid_i,
    input  logic       calc_i,
    input  logic       mode_i,
    input  logic       clear_i,

    output logic [4:0] result_o,
    output logic       output_valid_o
    );

    // add your implementation here

endmodule
